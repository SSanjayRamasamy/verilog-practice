module NAND_gate(input a,b,output y);
nand na1 (y,a,b);
endmodule