module NOR_gate(input a,b,y);
nor no1 (y,a,b);
endmodule