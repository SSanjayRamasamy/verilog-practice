module Barrel_Shifter #(parameter N=8)(input [N-1:0]data_in,input [$clog2(N)+1:0]shift,input [2:0]op,output [N-1:0]data_out);

endmodule