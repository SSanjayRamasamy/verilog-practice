module AND_gate (input a,b,output y);
and a1 (y,a,b);
endmodule