module XNOR_gate (input a,b,output y);
xnor xn1 (y,a,b);
endmodule