module Barrel_Shifter_tb();

endmodule